module LFSR_TB ();

    reg clk;
    reg rst;
    wire LFSR_out;

endmodule