// This is the top-level module that connects everything